module test;

    initial begin
        $display("hello world");
        $finish;
    end

endmodule