module test(input clock, input reset);

    initial begin
        $display("hello world");
        $finish;
    end

endmodule
