module relu(input clock, input reset);

    initial begin
        $display("hello from relu");
        $finish;
    end

endmodule
