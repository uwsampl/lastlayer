module adder(input clock, input reset);

    reg [31:0] r0;

endmodule
