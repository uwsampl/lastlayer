module __relu_dpi;


endmodule
