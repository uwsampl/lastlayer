module adder(input clock, input reset);

    initial begin
        $display("hello from adder");
        $finish;
    end

endmodule
