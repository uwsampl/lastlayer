module __adder_dpi;


endmodule
